LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
 
ENTITY add_8 IS
PORT ( a  : IN  std_logic_vector(7 DOWNTO 0);
       b  : IN  std_logic_vector(7 DOWNTO 0);
       s  : OUT std_logic_vector(7 DOWNTO 0) );
END add_8; 


